module TopModule(); 
	
	
endmodule