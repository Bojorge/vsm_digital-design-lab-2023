module VGA_controller ();




endmodule